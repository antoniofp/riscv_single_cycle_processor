module main(
	input clk
);
endmodule