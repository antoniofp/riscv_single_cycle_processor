module register_file (
	input clk, we3






);

endmodule